module and_gate(input x0, input x1, output y);
  assign y = x0 & x1;
endmodule

